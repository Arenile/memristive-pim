// Black Box
// black_box_1.v
// 
(* black_box *) module memristor (in, out);
inout in, out;
endmodule
